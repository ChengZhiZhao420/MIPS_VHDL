--Idenia Ayala
